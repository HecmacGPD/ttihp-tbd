magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771771680
<< checkpaint >>
rect -800 -1000 3680 63600
<< metal4 >>
rect 5922 62548 5982 62748
rect 6690 62548 6750 62748
rect 7458 62548 7518 62748
rect 8226 62548 8286 62748
rect 8994 62548 9054 62748
rect 9762 62548 9822 62748
rect 10530 62548 10590 62748
rect 11298 62548 11358 62748
rect 12066 62548 12126 62748
rect 12834 62548 12894 62748
rect 13602 62548 13662 62748
rect 14370 62548 14430 62748
rect 15138 62548 15198 62748
rect 15906 62548 15966 62748
rect 16674 62548 16734 62748
rect 17442 62548 17502 62748
rect 18210 62548 18270 62748
rect 18978 62548 19038 62748
rect 19746 62548 19806 62748
rect 20514 62548 20574 62748
rect 21282 62548 21342 62748
rect 22050 62548 22110 62748
rect 22818 62548 22878 62748
rect 23586 62548 23646 62748
rect 24354 62548 24414 62748
rect 25122 62548 25182 62748
rect 25890 62548 25950 62748
rect 26658 62548 26718 62748
rect 27426 62548 27486 62748
rect 28194 62548 28254 62748
rect 28962 62548 29022 62748
rect 29730 62548 29790 62748
rect 30498 62548 30558 62748
rect 31266 62548 31326 62748
rect 32034 62548 32094 62748
rect 32802 62548 32862 62748
rect 33570 62548 33630 62748
rect 34338 62548 34398 62748
rect 35106 62548 35166 62748
rect 35874 62548 35934 62748
rect 36642 62548 36702 62748
rect 37410 62548 37470 62748
rect 38178 62548 38238 62748
<< metal6 >>
rect 200 1000 680 61600
rect 1200 1000 1680 61600
rect 3761 0 4111 400
rect 8657 0 9007 400
rect 13553 0 13903 400
rect 18449 0 18799 400
rect 23345 0 23695 400
rect 28241 0 28591 400
rect 33137 0 33487 400
rect 38033 0 38383 400
<< labels >>
flabel metal4 s 37410 62548 37470 62748 0 FreeSans 320 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 38178 62548 38238 62748 0 FreeSans 320 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 36642 62548 36702 62748 0 FreeSans 320 90 0 0 rst_n
port 2 nsew signal input
flabel metal6 s 38033 0 38383 400 0 FreeSans 2624 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal6 s 33137 0 33487 400 0 FreeSans 2624 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal6 s 28241 0 28591 400 0 FreeSans 2624 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal6 s 23345 0 23695 400 0 FreeSans 2624 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal6 s 18449 0 18799 400 0 FreeSans 2624 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal6 s 13553 0 13903 400 0 FreeSans 2624 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal6 s 8657 0 9007 400 0 FreeSans 2624 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal6 s 3761 0 4111 400 0 FreeSans 2624 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 35874 62548 35934 62748 0 FreeSans 320 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 35106 62548 35166 62748 0 FreeSans 320 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 34338 62548 34398 62748 0 FreeSans 320 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 33570 62548 33630 62748 0 FreeSans 320 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 32802 62548 32862 62748 0 FreeSans 320 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 32034 62548 32094 62748 0 FreeSans 320 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 31266 62548 31326 62748 0 FreeSans 320 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 30498 62548 30558 62748 0 FreeSans 320 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 29730 62548 29790 62748 0 FreeSans 320 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 28962 62548 29022 62748 0 FreeSans 320 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 28194 62548 28254 62748 0 FreeSans 320 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 27426 62548 27486 62748 0 FreeSans 320 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 26658 62548 26718 62748 0 FreeSans 320 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 25890 62548 25950 62748 0 FreeSans 320 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 25122 62548 25182 62748 0 FreeSans 320 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 24354 62548 24414 62748 0 FreeSans 320 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 11298 62548 11358 62748 0 FreeSans 320 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 10530 62548 10590 62748 0 FreeSans 320 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 9762 62548 9822 62748 0 FreeSans 320 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8994 62548 9054 62748 0 FreeSans 320 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8226 62548 8286 62748 0 FreeSans 320 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7458 62548 7518 62748 0 FreeSans 320 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6690 62548 6750 62748 0 FreeSans 320 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 5922 62548 5982 62748 0 FreeSans 320 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 17442 62548 17502 62748 0 FreeSans 320 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 16674 62548 16734 62748 0 FreeSans 320 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 15906 62548 15966 62748 0 FreeSans 320 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 15138 62548 15198 62748 0 FreeSans 320 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 14370 62548 14430 62748 0 FreeSans 320 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 13602 62548 13662 62748 0 FreeSans 320 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12834 62548 12894 62748 0 FreeSans 320 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 12066 62548 12126 62748 0 FreeSans 320 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 23586 62548 23646 62748 0 FreeSans 320 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 22818 62548 22878 62748 0 FreeSans 320 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 22050 62548 22110 62748 0 FreeSans 320 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 21282 62548 21342 62748 0 FreeSans 320 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 20514 62548 20574 62748 0 FreeSans 320 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 19746 62548 19806 62748 0 FreeSans 320 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 18978 62548 19038 62748 0 FreeSans 320 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 18210 62548 18270 62748 0 FreeSans 320 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal6 200 1000 680 61600 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal6 1200 1000 1680 61600 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40416 62748
<< end >>
